 /*                                                                      
 Copyright 2020 Blue Liang, liangkangnan@163.com
                                                                         
 Licensed under the Apache License, Version 2.0 (the "License");         
 you may not use this file except in compliance with the License.        
 You may obtain a copy of the License at                                 
                                                                         
     http://www.apache.org/licenses/LICENSE-2.0                          
                                                                         
 Unless required by applicable law or agreed to in writing, software    
 distributed under the License is distributed on an "AS IS" BASIS,       
 WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 See the License for the specific language governing permissions and     
 limitations under the License.                                          
 */

`include "../core/defines.v"


module rom #(
    parameter DP = 4096)(

    input wire clk,
    input wire rst_n,
    input wire[31:0] addr_i,
    input wire[31:0] data_i,
    input wire[3:0] sel_i,
    input wire we_i,
	output wire[31:0] data_o,

    input wire req_valid_i,
    output wire req_ready_o,
    output wire rsp_valid_o,
    input wire rsp_ready_i
    );
wire[31:0] addr = addr_i[31:2];
//
//    gen_ram #(
//        .DP(DP),
//        .DW(32),
//        .MW(4),
//        .AW(32)
//    ) u_gen_ram(
//        .clk(clk),
//        .addr_i(addr),
//        .data_i(data_i),
//        .sel_i(sel_i),
//        .we_i(we_i),
//        .data_o(data_o)
//    );
wire [13:0] addr1;
assign addr1 = addr[13:0] ;
ram1 rom111 (
  .wr_data(data_i),    // input [31:0]
  .addr(addr1),          // input [13:0]
  .wr_en(we_i),        // input
  .clk(clk),            // input
  .rst(~rst_n),            // input
  .rd_data(data_o),     // output [31:0]
  .wr_byte_en(sel_i)
);

    vld_rdy #(
        .CUT_READY(0)
    ) u_vld_rdy(
        .clk(clk),
        .rst_n(rst_n),
        .vld_i(req_valid_i),
        .rdy_o(req_ready_o),
        .rdy_i(rsp_ready_i),
        .vld_o(rsp_valid_o)
    );

endmodule
